module fsm(e,w,clk,out)
output z;
input e, w, clk;
endmodule
